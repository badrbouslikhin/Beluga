.SUBCKT LM2731_33_BOOST_BLOCK_D1_WB_DIODE_ENCR A K
.include pspice://../LM2731_33_BOOST_BLOCK.D1.WB_DIODE.enl
XCALL A K LM2731_33_BOOST_BLOCK_D1_WB_DIODE 
.ENDS
