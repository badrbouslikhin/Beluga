***********************************
*     Created by WB Importer      *
***********************************
.SUBCKT LM2731_33_BOOST_BLOCK_Cout_WB_CAP_CERAMIC 2 4
*FAMILY = ANALOG
*FAMILY = ANALOG
R1 2 3 0.003
C1 3 4 4.698048442906574E-6 IC=0.0
R3 5 4 5; free space reduced by sqrt(dielectric constant)
R2 2 4 2.1285433987166873E8
R4 3 26 666666.6666666667
R6 3 7 666.6666666666667
C5 7 1 1.409414532871972E-7 IC=0.0
R7 3 10 66.66666666666669
C6 10 1 1.409414532871972E-7 IC=0.0
R8 3 13 6.666666666666668
C7 13 1 1.409414532871972E-7 IC=0.0
C2 26 1 1.409414532871972E-7 IC=0.0
R9 3 28 66666.66666666667
C3 28 1 1.409414532871972E-7 IC=0.0
R10 3 29 6666.666666666668
C4 29 1 1.409414532871972E-7 IC=0.0
L8 1 5 15p
R24 1 5 0.009000000000000001
L12 5 4 1n
.ENDS
