***********************************
*     Created by WB Importer      *
***********************************
.SUBCKT LM2731_33_BOOST_BLOCK_Cin_WB_CAP_POLARIZED 1 2
* C = 2.2E-6 F
* ESR = 0.0049 Ohm

Ccap 1 3 2.2E-6
Resr 3 2 0.0049

.ENDS
