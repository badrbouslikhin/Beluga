***********************************
*     Created by WB Importer      *
***********************************
.subckt LM2731_33_BOOST_BLOCK_WB_LM27313_BOOST_BLOCK_Rp 1 2
Rp 1 2 51000.0

.ends
