***********************************
*     Created by WB Importer      *
***********************************
.subckt LM2731_33_BOOST_BLOCK_WB_LM27313_BOOST_BLOCK_Cf 6 5
Cf 6 5 1.0E-10

.ends
