***********************************
*     Created by WB Importer      *
***********************************
.SUBCKT INPUT_BLOCK_Vin_WB_STARTUP_VOLTAGE_SOURCE 1 2
Rsource 3 1 1m
Vin1 3 2 PULSE 0 5.0 1u 1m
.ENDS
