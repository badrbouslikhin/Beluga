***********************************
*     Created by WB Importer      *
***********************************
.subckt LM2731_33_BOOST_BLOCK_WB_LM27313_BOOST_BLOCK_Rfbb 5 0
Rfbb 5 0 13300.0

.ends
